
//================================================================================================
// Version  Date         Who  What
//----------------------------------------------------------------------
//   1.0.0  08-Jun-2025  DWW  Initial creation
//================================================================================================
localparam RTL_TYPE      = 52125;
localparam RTL_SUBTYPE   = 0;

localparam VERSION_MAJOR = 1;
localparam VERSION_MINOR = 0;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 0;

